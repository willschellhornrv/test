module rom_file(out, address);

	// 2^10 inputs, so 1024 indices
	input [9:0] address;
	output out;
	reg out;
	
 always @ (address) begin
	case (address)
		0 : out = 1'b0;
		1 : out = 1'b0;
		2 : out = 1'b1;
		3 : out = 1'b1;
		4 : out = 1'b0;
		5 : out = 1'b1;
		6 : out = 1'b0;
		7 : out = 1'b1;
		8 : out = 1'b0;
		9 : out = 1'b0;
		10 : out = 1'b0;
		11 : out = 1'b1;
		12 : out = 1'b0;
		13 : out = 1'b1;
		14 : out = 1'b0;
		15 : out = 1'b0;
		16 : out = 1'b0;
		17 : out = 1'b1;
		18 : out = 1'b0;
		19 : out = 1'b1;
		20 : out = 1'b0;
		21 : out = 1'b0;
		22 : out = 1'b0;
		23 : out = 1'b1;
		24 : out = 1'b0;
		25 : out = 1'b0;
		26 : out = 1'b0;
		27 : out = 1'b0;
		28 : out = 1'b0;
		29 : out = 1'b1;
		30 : out = 1'b0;
		31 : out = 1'b1;
		32 : out = 1'b0;
		33 : out = 1'b0;
		34 : out = 1'b0;
		35 : out = 1'b0;
		36 : out = 1'b0;
		37 : out = 1'b1;
		38 : out = 1'b0;
		39 : out = 1'b0;
		40 : out = 1'b0;
		41 : out = 1'b1;
		42 : out = 1'b0;
		43 : out = 1'b1;
		44 : out = 1'b0;
		45 : out = 1'b0;
		46 : out = 1'b0;
		47 : out = 1'b1;
		48 : out = 1'b0;
		49 : out = 1'b0;
		50 : out = 1'b0;
		51 : out = 1'b0;
		52 : out = 1'b0;
		53 : out = 1'b1;
		54 : out = 1'b0;
		55 : out = 1'b0;
		56 : out = 1'b0;
		57 : out = 1'b0;
		58 : out = 1'b0;
		59 : out = 1'b1;
		60 : out = 1'b0;
		61 : out = 1'b1;
		62 : out = 1'b0;
		63 : out = 1'b0;
		64 : out = 1'b0;
		65 : out = 1'b0;
		66 : out = 1'b0;
		67 : out = 1'b1;
		68 : out = 1'b0;
		69 : out = 1'b0;
		70 : out = 1'b0;
		71 : out = 1'b1;
		72 : out = 1'b0;
		73 : out = 1'b1;
		74 : out = 1'b0;
		75 : out = 1'b0;
		76 : out = 1'b0;
		77 : out = 1'b0;
		78 : out = 1'b0;
		79 : out = 1'b1;
		80 : out = 1'b0;
		81 : out = 1'b0;
		82 : out = 1'b0;
		83 : out = 1'b1;
		84 : out = 1'b0;
		85 : out = 1'b0;
		86 : out = 1'b0;
		87 : out = 1'b0;
		88 : out = 1'b0;
		89 : out = 1'b1;
		90 : out = 1'b0;
		91 : out = 1'b0;
		92 : out = 1'b0;
		93 : out = 1'b0;
		94 : out = 1'b0;
		95 : out = 1'b0;
		96 : out = 1'b0;
		97 : out = 1'b1;
		98 : out = 1'b0;
		99 : out = 1'b0;
		100 : out = 1'b0;
		101 : out = 1'b1;
		102 : out = 1'b0;
		103 : out = 1'b1;
		104 : out = 1'b0;
		105 : out = 1'b0;
		106 : out = 1'b0;
		107 : out = 1'b1;
		108 : out = 1'b0;
		109 : out = 1'b1;
		110 : out = 1'b0;
		111 : out = 1'b0;
		112 : out = 1'b0;
		113 : out = 1'b1;
		114 : out = 1'b0;
		115 : out = 1'b0;
		116 : out = 1'b0;
		117 : out = 1'b0;
		118 : out = 1'b0;
		119 : out = 1'b0;
		120 : out = 1'b0;
		121 : out = 1'b0;
		122 : out = 1'b0;
		123 : out = 1'b0;
		124 : out = 1'b0;
		125 : out = 1'b0;
		126 : out = 1'b0;
		127 : out = 1'b1;
		128 : out = 1'b0;
		129 : out = 1'b0;
		130 : out = 1'b0;
		131 : out = 1'b1;
		132 : out = 1'b0;
		133 : out = 1'b0;
		134 : out = 1'b0;
		135 : out = 1'b0;
		136 : out = 1'b0;
		137 : out = 1'b1;
		138 : out = 1'b0;
		139 : out = 1'b1;
		140 : out = 1'b0;
		141 : out = 1'b0;
		142 : out = 1'b0;
		143 : out = 1'b0;
		144 : out = 1'b0;
		145 : out = 1'b0;
		146 : out = 1'b0;
		147 : out = 1'b0;
		148 : out = 1'b0;
		149 : out = 1'b1;
		150 : out = 1'b0;
		151 : out = 1'b1;
		152 : out = 1'b0;
		153 : out = 1'b0;
		154 : out = 1'b0;
		155 : out = 1'b0;
		156 : out = 1'b0;
		157 : out = 1'b1;
		158 : out = 1'b0;
		159 : out = 1'b0;
		160 : out = 1'b0;
		161 : out = 1'b0;
		162 : out = 1'b0;
		163 : out = 1'b1;
		164 : out = 1'b0;
		165 : out = 1'b0;
		166 : out = 1'b0;
		167 : out = 1'b1;
		168 : out = 1'b0;
		169 : out = 1'b0;
		170 : out = 1'b0;
		171 : out = 1'b0;
		172 : out = 1'b0;
		173 : out = 1'b1;
		174 : out = 1'b0;
		175 : out = 1'b0;
		176 : out = 1'b0;
		177 : out = 1'b0;
		178 : out = 1'b0;
		179 : out = 1'b1;
		180 : out = 1'b0;
		181 : out = 1'b1;
		182 : out = 1'b0;
		183 : out = 1'b0;
		184 : out = 1'b0;
		185 : out = 1'b0;
		186 : out = 1'b0;
		187 : out = 1'b0;
		188 : out = 1'b0;
		189 : out = 1'b0;
		190 : out = 1'b0;
		191 : out = 1'b1;
		192 : out = 1'b0;
		193 : out = 1'b1;
		194 : out = 1'b0;
		195 : out = 1'b0;
		196 : out = 1'b0;
		197 : out = 1'b1;
		198 : out = 1'b0;
		199 : out = 1'b1;
		200 : out = 1'b0;
		201 : out = 1'b0;
		202 : out = 1'b0;
		203 : out = 1'b0;
		204 : out = 1'b0;
		205 : out = 1'b0;
		206 : out = 1'b0;
		207 : out = 1'b0;
		208 : out = 1'b0;
		209 : out = 1'b0;
		210 : out = 1'b0;
		211 : out = 1'b1;
		212 : out = 1'b0;
		213 : out = 1'b0;
		214 : out = 1'b0;
		215 : out = 1'b0;
		216 : out = 1'b0;
		217 : out = 1'b0;
		218 : out = 1'b0;
		219 : out = 1'b0;
		220 : out = 1'b0;
		221 : out = 1'b0;
		222 : out = 1'b0;
		223 : out = 1'b1;
		224 : out = 1'b0;
		225 : out = 1'b0;
		226 : out = 1'b0;
		227 : out = 1'b1;
		228 : out = 1'b0;
		229 : out = 1'b1;
		230 : out = 1'b0;
		231 : out = 1'b0;
		232 : out = 1'b0;
		233 : out = 1'b1;
		234 : out = 1'b0;
		235 : out = 1'b0;
		236 : out = 1'b0;
		237 : out = 1'b0;
		238 : out = 1'b0;
		239 : out = 1'b1;
		240 : out = 1'b0;
		241 : out = 1'b1;
		242 : out = 1'b0;
		243 : out = 1'b0;
		244 : out = 1'b0;
		245 : out = 1'b0;
		246 : out = 1'b0;
		247 : out = 1'b0;
		248 : out = 1'b0;
		249 : out = 1'b0;
		250 : out = 1'b0;
		251 : out = 1'b1;
		252 : out = 1'b0;
		253 : out = 1'b0;
		254 : out = 1'b0;
		255 : out = 1'b0;
		256 : out = 1'b0;
		257 : out = 1'b1;
		258 : out = 1'b0;
		259 : out = 1'b0;
		260 : out = 1'b0;
		261 : out = 1'b0;
		262 : out = 1'b0;
		263 : out = 1'b1;
		264 : out = 1'b0;
		265 : out = 1'b0;
		266 : out = 1'b0;
		267 : out = 1'b0;
		268 : out = 1'b0;
		269 : out = 1'b1;
		270 : out = 1'b0;
		271 : out = 1'b1;
		272 : out = 1'b0;
		273 : out = 1'b0;
		274 : out = 1'b0;
		275 : out = 1'b0;
		276 : out = 1'b0;
		277 : out = 1'b1;
		278 : out = 1'b0;
		279 : out = 1'b0;
		280 : out = 1'b0;
		281 : out = 1'b1;
		282 : out = 1'b0;
		283 : out = 1'b1;
		284 : out = 1'b0;
		285 : out = 1'b0;
		286 : out = 1'b0;
		287 : out = 1'b0;
		288 : out = 1'b0;
		289 : out = 1'b0;
		290 : out = 1'b0;
		291 : out = 1'b0;
		292 : out = 1'b0;
		293 : out = 1'b1;
		294 : out = 1'b0;
		295 : out = 1'b0;
		296 : out = 1'b0;
		297 : out = 1'b0;
		298 : out = 1'b0;
		299 : out = 1'b0;
		300 : out = 1'b0;
		301 : out = 1'b0;
		302 : out = 1'b0;
		303 : out = 1'b0;
		304 : out = 1'b0;
		305 : out = 1'b0;
		306 : out = 1'b0;
		307 : out = 1'b1;
		308 : out = 1'b0;
		309 : out = 1'b0;
		310 : out = 1'b0;
		311 : out = 1'b1;
		312 : out = 1'b0;
		313 : out = 1'b1;
		314 : out = 1'b0;
		315 : out = 1'b0;
		316 : out = 1'b0;
		317 : out = 1'b1;
		318 : out = 1'b0;
		319 : out = 1'b0;
		320 : out = 1'b0;
		321 : out = 1'b0;
		322 : out = 1'b0;
		323 : out = 1'b0;
		324 : out = 1'b0;
		325 : out = 1'b0;
		326 : out = 1'b0;
		327 : out = 1'b0;
		328 : out = 1'b0;
		329 : out = 1'b0;
		330 : out = 1'b0;
		331 : out = 1'b1;
		332 : out = 1'b0;
		333 : out = 1'b0;
		334 : out = 1'b0;
		335 : out = 1'b0;
		336 : out = 1'b0;
		337 : out = 1'b1;
		338 : out = 1'b0;
		339 : out = 1'b0;
		340 : out = 1'b0;
		341 : out = 1'b0;
		342 : out = 1'b0;
		343 : out = 1'b0;
		344 : out = 1'b0;
		345 : out = 1'b0;
		346 : out = 1'b0;
		347 : out = 1'b1;
		348 : out = 1'b0;
		349 : out = 1'b1;
		350 : out = 1'b0;
		351 : out = 1'b0;
		352 : out = 1'b0;
		353 : out = 1'b1;
		354 : out = 1'b0;
		355 : out = 1'b0;
		356 : out = 1'b0;
		357 : out = 1'b0;
		358 : out = 1'b0;
		359 : out = 1'b1;
		360 : out = 1'b0;
		361 : out = 1'b0;
		362 : out = 1'b0;
		363 : out = 1'b0;
		364 : out = 1'b0;
		365 : out = 1'b0;
		366 : out = 1'b0;
		367 : out = 1'b1;
		368 : out = 1'b0;
		369 : out = 1'b0;
		370 : out = 1'b0;
		371 : out = 1'b0;
		372 : out = 1'b0;
		373 : out = 1'b1;
		374 : out = 1'b0;
		375 : out = 1'b0;
		376 : out = 1'b0;
		377 : out = 1'b0;
		378 : out = 1'b0;
		379 : out = 1'b1;
		380 : out = 1'b0;
		381 : out = 1'b0;
		382 : out = 1'b0;
		383 : out = 1'b1;
		384 : out = 1'b0;
		385 : out = 1'b0;
		386 : out = 1'b0;
		387 : out = 1'b0;
		388 : out = 1'b0;
		389 : out = 1'b1;
		390 : out = 1'b0;
		391 : out = 1'b0;
		392 : out = 1'b0;
		393 : out = 1'b0;
		394 : out = 1'b0;
		395 : out = 1'b0;
		396 : out = 1'b0;
		397 : out = 1'b1;
		398 : out = 1'b0;
		399 : out = 1'b0;
		400 : out = 1'b0;
		401 : out = 1'b1;
		402 : out = 1'b0;
		403 : out = 1'b0;
		404 : out = 1'b0;
		405 : out = 1'b0;
		406 : out = 1'b0;
		407 : out = 1'b0;
		408 : out = 1'b0;
		409 : out = 1'b1;
		410 : out = 1'b0;
		411 : out = 1'b0;
		412 : out = 1'b0;
		413 : out = 1'b0;
		414 : out = 1'b0;
		415 : out = 1'b0;
		416 : out = 1'b0;
		417 : out = 1'b0;
		418 : out = 1'b0;
		419 : out = 1'b1;
		420 : out = 1'b0;
		421 : out = 1'b1;
		422 : out = 1'b0;
		423 : out = 1'b0;
		424 : out = 1'b0;
		425 : out = 1'b0;
		426 : out = 1'b0;
		427 : out = 1'b0;
		428 : out = 1'b0;
		429 : out = 1'b0;
		430 : out = 1'b0;
		431 : out = 1'b1;
		432 : out = 1'b0;
		433 : out = 1'b1;
		434 : out = 1'b0;
		435 : out = 1'b0;
		436 : out = 1'b0;
		437 : out = 1'b0;
		438 : out = 1'b0;
		439 : out = 1'b1;
		440 : out = 1'b0;
		441 : out = 1'b0;
		442 : out = 1'b0;
		443 : out = 1'b1;
		444 : out = 1'b0;
		445 : out = 1'b0;
		446 : out = 1'b0;
		447 : out = 1'b0;
		448 : out = 1'b0;
		449 : out = 1'b1;
		450 : out = 1'b0;
		451 : out = 1'b0;
		452 : out = 1'b0;
		453 : out = 1'b0;
		454 : out = 1'b0;
		455 : out = 1'b0;
		456 : out = 1'b0;
		457 : out = 1'b1;
		458 : out = 1'b0;
		459 : out = 1'b0;
		460 : out = 1'b0;
		461 : out = 1'b1;
		462 : out = 1'b0;
		463 : out = 1'b1;
		464 : out = 1'b0;
		465 : out = 1'b0;
		466 : out = 1'b0;
		467 : out = 1'b1;
		468 : out = 1'b0;
		469 : out = 1'b0;
		470 : out = 1'b0;
		471 : out = 1'b0;
		472 : out = 1'b0;
		473 : out = 1'b0;
		474 : out = 1'b0;
		475 : out = 1'b0;
		476 : out = 1'b0;
		477 : out = 1'b0;
		478 : out = 1'b0;
		479 : out = 1'b1;
		480 : out = 1'b0;
		481 : out = 1'b0;
		482 : out = 1'b0;
		483 : out = 1'b0;
		484 : out = 1'b0;
		485 : out = 1'b0;
		486 : out = 1'b0;
		487 : out = 1'b1;
		488 : out = 1'b0;
		489 : out = 1'b0;
		490 : out = 1'b0;
		491 : out = 1'b1;
		492 : out = 1'b0;
		493 : out = 1'b0;
		494 : out = 1'b0;
		495 : out = 1'b0;
		496 : out = 1'b0;
		497 : out = 1'b0;
		498 : out = 1'b0;
		499 : out = 1'b1;
		500 : out = 1'b0;
		501 : out = 1'b0;
		502 : out = 1'b0;
		503 : out = 1'b1;
		504 : out = 1'b0;
		505 : out = 1'b0;
		506 : out = 1'b0;
		507 : out = 1'b0;
		508 : out = 1'b0;
		509 : out = 1'b1;
		510 : out = 1'b0;
		511 : out = 1'b0;
		512 : out = 1'b0;
		513 : out = 1'b0;
		514 : out = 1'b0;
		515 : out = 1'b0;
		516 : out = 1'b0;
		517 : out = 1'b0;
		518 : out = 1'b0;
		519 : out = 1'b0;
		520 : out = 1'b0;
		521 : out = 1'b1;
		522 : out = 1'b0;
		523 : out = 1'b1;
		524 : out = 1'b0;
		525 : out = 1'b0;
		526 : out = 1'b0;
		527 : out = 1'b0;
		528 : out = 1'b0;
		529 : out = 1'b0;
		530 : out = 1'b0;
		531 : out = 1'b0;
		532 : out = 1'b0;
		533 : out = 1'b0;
		534 : out = 1'b0;
		535 : out = 1'b0;
		536 : out = 1'b0;
		537 : out = 1'b0;
		538 : out = 1'b0;
		539 : out = 1'b0;
		540 : out = 1'b0;
		541 : out = 1'b1;
		542 : out = 1'b0;
		543 : out = 1'b0;
		544 : out = 1'b0;
		545 : out = 1'b0;
		546 : out = 1'b0;
		547 : out = 1'b1;
		548 : out = 1'b0;
		549 : out = 1'b0;
		550 : out = 1'b0;
		551 : out = 1'b0;
		552 : out = 1'b0;
		553 : out = 1'b0;
		554 : out = 1'b0;
		555 : out = 1'b0;
		556 : out = 1'b0;
		557 : out = 1'b1;
		558 : out = 1'b0;
		559 : out = 1'b0;
		560 : out = 1'b0;
		561 : out = 1'b0;
		562 : out = 1'b0;
		563 : out = 1'b1;
		564 : out = 1'b0;
		565 : out = 1'b0;
		566 : out = 1'b0;
		567 : out = 1'b0;
		568 : out = 1'b0;
		569 : out = 1'b1;
		570 : out = 1'b0;
		571 : out = 1'b1;
		572 : out = 1'b0;
		573 : out = 1'b0;
		574 : out = 1'b0;
		575 : out = 1'b0;
		576 : out = 1'b0;
		577 : out = 1'b1;
		578 : out = 1'b0;
		579 : out = 1'b0;
		580 : out = 1'b0;
		581 : out = 1'b0;
		582 : out = 1'b0;
		583 : out = 1'b0;
		584 : out = 1'b0;
		585 : out = 1'b0;
		586 : out = 1'b0;
		587 : out = 1'b1;
		588 : out = 1'b0;
		589 : out = 1'b0;
		590 : out = 1'b0;
		591 : out = 1'b0;
		592 : out = 1'b0;
		593 : out = 1'b1;
		594 : out = 1'b0;
		595 : out = 1'b0;
		596 : out = 1'b0;
		597 : out = 1'b0;
		598 : out = 1'b0;
		599 : out = 1'b1;
		600 : out = 1'b0;
		601 : out = 1'b1;
		602 : out = 1'b0;
		603 : out = 1'b0;
		604 : out = 1'b0;
		605 : out = 1'b0;
		606 : out = 1'b0;
		607 : out = 1'b1;
		608 : out = 1'b0;
		609 : out = 1'b0;
		610 : out = 1'b0;
		611 : out = 1'b0;
		612 : out = 1'b0;
		613 : out = 1'b1;
		614 : out = 1'b0;
		615 : out = 1'b0;
		616 : out = 1'b0;
		617 : out = 1'b1;
		618 : out = 1'b0;
		619 : out = 1'b1;
		620 : out = 1'b0;
		621 : out = 1'b0;
		622 : out = 1'b0;
		623 : out = 1'b0;
		624 : out = 1'b0;
		625 : out = 1'b0;
		626 : out = 1'b0;
		627 : out = 1'b0;
		628 : out = 1'b0;
		629 : out = 1'b0;
		630 : out = 1'b0;
		631 : out = 1'b1;
		632 : out = 1'b0;
		633 : out = 1'b0;
		634 : out = 1'b0;
		635 : out = 1'b0;
		636 : out = 1'b0;
		637 : out = 1'b0;
		638 : out = 1'b0;
		639 : out = 1'b0;
		640 : out = 1'b0;
		641 : out = 1'b1;
		642 : out = 1'b0;
		643 : out = 1'b1;
		644 : out = 1'b0;
		645 : out = 1'b0;
		646 : out = 1'b0;
		647 : out = 1'b1;
		648 : out = 1'b0;
		649 : out = 1'b0;
		650 : out = 1'b0;
		651 : out = 1'b0;
		652 : out = 1'b0;
		653 : out = 1'b1;
		654 : out = 1'b0;
		655 : out = 1'b0;
		656 : out = 1'b0;
		657 : out = 1'b0;
		658 : out = 1'b0;
		659 : out = 1'b1;
		660 : out = 1'b0;
		661 : out = 1'b1;
		662 : out = 1'b0;
		663 : out = 1'b0;
		664 : out = 1'b0;
		665 : out = 1'b0;
		666 : out = 1'b0;
		667 : out = 1'b0;
		668 : out = 1'b0;
		669 : out = 1'b0;
		670 : out = 1'b0;
		671 : out = 1'b0;
		672 : out = 1'b0;
		673 : out = 1'b1;
		674 : out = 1'b0;
		675 : out = 1'b0;
		676 : out = 1'b0;
		677 : out = 1'b1;
		678 : out = 1'b0;
		679 : out = 1'b0;
		680 : out = 1'b0;
		681 : out = 1'b0;
		682 : out = 1'b0;
		683 : out = 1'b1;
		684 : out = 1'b0;
		685 : out = 1'b0;
		686 : out = 1'b0;
		687 : out = 1'b0;
		688 : out = 1'b0;
		689 : out = 1'b0;
		690 : out = 1'b0;
		691 : out = 1'b1;
		692 : out = 1'b0;
		693 : out = 1'b0;
		694 : out = 1'b0;
		695 : out = 1'b0;
		696 : out = 1'b0;
		697 : out = 1'b0;
		698 : out = 1'b0;
		699 : out = 1'b0;
		700 : out = 1'b0;
		701 : out = 1'b1;
		702 : out = 1'b0;
		703 : out = 1'b0;
		704 : out = 1'b0;
		705 : out = 1'b0;
		706 : out = 1'b0;
		707 : out = 1'b0;
		708 : out = 1'b0;
		709 : out = 1'b1;
		710 : out = 1'b0;
		711 : out = 1'b0;
		712 : out = 1'b0;
		713 : out = 1'b0;
		714 : out = 1'b0;
		715 : out = 1'b0;
		716 : out = 1'b0;
		717 : out = 1'b0;
		718 : out = 1'b0;
		719 : out = 1'b1;
		720 : out = 1'b0;
		721 : out = 1'b0;
		722 : out = 1'b0;
		723 : out = 1'b0;
		724 : out = 1'b0;
		725 : out = 1'b0;
		726 : out = 1'b0;
		727 : out = 1'b1;
		728 : out = 1'b0;
		729 : out = 1'b0;
		730 : out = 1'b0;
		731 : out = 1'b0;
		732 : out = 1'b0;
		733 : out = 1'b1;
		734 : out = 1'b0;
		735 : out = 1'b0;
		736 : out = 1'b0;
		737 : out = 1'b0;
		738 : out = 1'b0;
		739 : out = 1'b1;
		740 : out = 1'b0;
		741 : out = 1'b0;
		742 : out = 1'b0;
		743 : out = 1'b1;
		744 : out = 1'b0;
		745 : out = 1'b0;
		746 : out = 1'b0;
		747 : out = 1'b0;
		748 : out = 1'b0;
		749 : out = 1'b0;
		750 : out = 1'b0;
		751 : out = 1'b1;
		752 : out = 1'b0;
		753 : out = 1'b0;
		754 : out = 1'b0;
		755 : out = 1'b0;
		756 : out = 1'b0;
		757 : out = 1'b1;
		758 : out = 1'b0;
		759 : out = 1'b0;
		760 : out = 1'b0;
		761 : out = 1'b1;
		762 : out = 1'b0;
		763 : out = 1'b0;
		764 : out = 1'b0;
		765 : out = 1'b0;
		766 : out = 1'b0;
		767 : out = 1'b0;
		768 : out = 1'b0;
		769 : out = 1'b1;
		770 : out = 1'b0;
		771 : out = 1'b0;
		772 : out = 1'b0;
		773 : out = 1'b1;
		774 : out = 1'b0;
		775 : out = 1'b0;
		776 : out = 1'b0;
		777 : out = 1'b0;
		778 : out = 1'b0;
		779 : out = 1'b0;
		780 : out = 1'b0;
		781 : out = 1'b0;
		782 : out = 1'b0;
		783 : out = 1'b0;
		784 : out = 1'b0;
		785 : out = 1'b0;
		786 : out = 1'b0;
		787 : out = 1'b1;
		788 : out = 1'b0;
		789 : out = 1'b0;
		790 : out = 1'b0;
		791 : out = 1'b0;
		792 : out = 1'b0;
		793 : out = 1'b0;
		794 : out = 1'b0;
		795 : out = 1'b0;
		796 : out = 1'b0;
		797 : out = 1'b1;
		798 : out = 1'b0;
		799 : out = 1'b0;
		800 : out = 1'b0;
		801 : out = 1'b0;
		802 : out = 1'b0;
		803 : out = 1'b0;
		804 : out = 1'b0;
		805 : out = 1'b0;
		806 : out = 1'b0;
		807 : out = 1'b0;
		808 : out = 1'b0;
		809 : out = 1'b1;
		810 : out = 1'b0;
		811 : out = 1'b1;
		812 : out = 1'b0;
		813 : out = 1'b0;
		814 : out = 1'b0;
		815 : out = 1'b0;
		816 : out = 1'b0;
		817 : out = 1'b0;
		818 : out = 1'b0;
		819 : out = 1'b0;
		820 : out = 1'b0;
		821 : out = 1'b1;
		822 : out = 1'b0;
		823 : out = 1'b1;
		824 : out = 1'b0;
		825 : out = 1'b0;
		826 : out = 1'b0;
		827 : out = 1'b1;
		828 : out = 1'b0;
		829 : out = 1'b1;
		830 : out = 1'b0;
		831 : out = 1'b0;
		832 : out = 1'b0;
		833 : out = 1'b0;
		834 : out = 1'b0;
		835 : out = 1'b0;
		836 : out = 1'b0;
		837 : out = 1'b0;
		838 : out = 1'b0;
		839 : out = 1'b1;
		840 : out = 1'b0;
		841 : out = 1'b0;
		842 : out = 1'b0;
		843 : out = 1'b0;
		844 : out = 1'b0;
		845 : out = 1'b0;
		846 : out = 1'b0;
		847 : out = 1'b0;
		848 : out = 1'b0;
		849 : out = 1'b0;
		850 : out = 1'b0;
		851 : out = 1'b0;
		852 : out = 1'b0;
		853 : out = 1'b1;
		854 : out = 1'b0;
		855 : out = 1'b0;
		856 : out = 1'b0;
		857 : out = 1'b1;
		858 : out = 1'b0;
		859 : out = 1'b1;
		860 : out = 1'b0;
		861 : out = 1'b0;
		862 : out = 1'b0;
		863 : out = 1'b1;
		864 : out = 1'b0;
		865 : out = 1'b0;
		866 : out = 1'b0;
		867 : out = 1'b0;
		868 : out = 1'b0;
		869 : out = 1'b0;
		870 : out = 1'b0;
		871 : out = 1'b0;
		872 : out = 1'b0;
		873 : out = 1'b0;
		874 : out = 1'b0;
		875 : out = 1'b0;
		876 : out = 1'b0;
		877 : out = 1'b1;
		878 : out = 1'b0;
		879 : out = 1'b0;
		880 : out = 1'b0;
		881 : out = 1'b1;
		882 : out = 1'b0;
		883 : out = 1'b1;
		884 : out = 1'b0;
		885 : out = 1'b0;
		886 : out = 1'b0;
		887 : out = 1'b1;
		888 : out = 1'b0;
		889 : out = 1'b0;
		890 : out = 1'b0;
		891 : out = 1'b0;
		892 : out = 1'b0;
		893 : out = 1'b0;
		894 : out = 1'b0;
		895 : out = 1'b0;
		896 : out = 1'b0;
		897 : out = 1'b0;
		898 : out = 1'b0;
		899 : out = 1'b0;
		900 : out = 1'b0;
		901 : out = 1'b0;
		902 : out = 1'b0;
		903 : out = 1'b0;
		904 : out = 1'b0;
		905 : out = 1'b0;
		906 : out = 1'b0;
		907 : out = 1'b1;
		908 : out = 1'b0;
		909 : out = 1'b0;
		910 : out = 1'b0;
		911 : out = 1'b1;
		912 : out = 1'b0;
		913 : out = 1'b0;
		914 : out = 1'b0;
		915 : out = 1'b0;
		916 : out = 1'b0;
		917 : out = 1'b0;
		918 : out = 1'b0;
		919 : out = 1'b1;
		920 : out = 1'b0;
		921 : out = 1'b0;
		922 : out = 1'b0;
		923 : out = 1'b0;
		924 : out = 1'b0;
		925 : out = 1'b0;
		926 : out = 1'b0;
		927 : out = 1'b0;
		928 : out = 1'b0;
		929 : out = 1'b1;
		930 : out = 1'b0;
		931 : out = 1'b0;
		932 : out = 1'b0;
		933 : out = 1'b0;
		934 : out = 1'b0;
		935 : out = 1'b0;
		936 : out = 1'b0;
		937 : out = 1'b1;
		938 : out = 1'b0;
		939 : out = 1'b0;
		940 : out = 1'b0;
		941 : out = 1'b1;
		942 : out = 1'b0;
		943 : out = 1'b0;
		944 : out = 1'b0;
		945 : out = 1'b0;
		946 : out = 1'b0;
		947 : out = 1'b1;
		948 : out = 1'b0;
		949 : out = 1'b0;
		950 : out = 1'b0;
		951 : out = 1'b0;
		952 : out = 1'b0;
		953 : out = 1'b1;
		954 : out = 1'b0;
		955 : out = 1'b0;
		956 : out = 1'b0;
		957 : out = 1'b0;
		958 : out = 1'b0;
		959 : out = 1'b0;
		960 : out = 1'b0;
		961 : out = 1'b0;
		962 : out = 1'b0;
		963 : out = 1'b0;
		964 : out = 1'b0;
		965 : out = 1'b0;
		966 : out = 1'b0;
		967 : out = 1'b1;
		968 : out = 1'b0;
		969 : out = 1'b0;
		970 : out = 1'b0;
		971 : out = 1'b1;
		972 : out = 1'b0;
		973 : out = 1'b0;
		974 : out = 1'b0;
		975 : out = 1'b0;
		976 : out = 1'b0;
		977 : out = 1'b1;
		978 : out = 1'b0;
		979 : out = 1'b0;
		980 : out = 1'b0;
		981 : out = 1'b0;
		982 : out = 1'b0;
		983 : out = 1'b1;
		984 : out = 1'b0;
		985 : out = 1'b0;
		986 : out = 1'b0;
		987 : out = 1'b0;
		988 : out = 1'b0;
		989 : out = 1'b0;
		990 : out = 1'b0;
		991 : out = 1'b1;
		992 : out = 1'b0;
		993 : out = 1'b0;
		994 : out = 1'b0;
		995 : out = 1'b0;
		996 : out = 1'b0;
		997 : out = 1'b1;
		998 : out = 1'b0;
		999 : out = 1'b0;
		1000 : out = 1'b0;
		1001 : out = 1'b0;
		1002 : out = 1'b0;
		1003 : out = 1'b0;
		1004 : out = 1'b0;
		1005 : out = 1'b0;
		1006 : out = 1'b0;
		1007 : out = 1'b0;
		1008 : out = 1'b0;
		1009 : out = 1'b1;
		1010 : out = 1'b0;
		1011 : out = 1'b0;
		1012 : out = 1'b0;
		1013 : out = 1'b1;
		1014 : out = 1'b0;
		1015 : out = 1'b0;
		1016 : out = 1'b0;
		1017 : out = 1'b0;
		1018 : out = 1'b0;
		1019 : out = 1'b1;
		1020 : out = 1'b0;
		1021 : out = 1'b1;
		1022 : out = 1'b0;
		1023 : out = 1'b0;
	endcase
end
		

endmodule
